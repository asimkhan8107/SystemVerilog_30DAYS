module design_block(output bit [7:0] addr);
  initial
    begin
      	addr <= 10;
    end
endmodule
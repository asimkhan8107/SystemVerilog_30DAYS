module adder(
  	input [3:0] a,b,
  	output [6:0] sum
	);
  
  assign sum = a + b;
endmodule
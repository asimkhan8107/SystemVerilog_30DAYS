/*				Array Callback				*/
`include "slave_driver.sv"
`include "slave_env.sv"
`include "error_test.sv"
interface intf;
  // declaring signals
  logic [3:0] a,b;
  logic [6:0] sum;
endinterface